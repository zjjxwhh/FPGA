library verilog;
use verilog.vl_types.all;
entity seg_driver_tb is
end seg_driver_tb;
