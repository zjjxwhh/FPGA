library verilog;
use verilog.vl_types.all;
entity top1_tb is
end top1_tb;
