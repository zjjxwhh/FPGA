`timescale 1ns/1ps
module top1_tb;

	reg a;
	reg b;
	reg c;
	
	wire d;

	top1 top1_inst(
		.a(a), 
		.b(b),
		.c(c), 
		.d(d)
	);
	
	initial
	begin
		a = 0; b = 0; c = 0;
		#200
		a = 0; b = 0; c = 1;
		#200
		a = 0; b = 1; c = 0;
		#200
		a = 0; b = 1; c = 1;
		#200
		a = 1; b = 0; c = 0;
		#200
		a = 1; b = 0; c = 1;
		#200
		a = 1; b = 1; c = 0;
		#200
		a = 1; b = 1; c = 1;
		#200
		$stop;
	end

endmodule 
