library verilog;
use verilog.vl_types.all;
entity and_gate_tb is
end and_gate_tb;
