library verilog;
use verilog.vl_types.all;
entity digital_clock_tb is
end digital_clock_tb;
