library verilog;
use verilog.vl_types.all;
entity led_driver_tb is
end led_driver_tb;
