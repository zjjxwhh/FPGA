library verilog;
use verilog.vl_types.all;
entity top1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : out    vl_logic
    );
end top1;
