library verilog;
use verilog.vl_types.all;
entity calculator_tb is
end calculator_tb;
